/*
    注意事项:
    rstn 表示 rst 取非
    当 block_l2 == 1 时, 所有寄存器保持原值
    当 rstn == 0 或 clear_l2 == 1 时, 所有寄存器清零
    其他情况 xxx_l2 = xxx_l1

*/


module L2 (
    input  wire        clk,
    input  wire        rstn,
    input  wire        clear_l2,
    input  wire        block_l2,
    input  wire [31:0] pc_l1,
    input  wire [31:0] imm_l1,
    input  wire [ 4:0] rd_l1,
    input  wire [ 4:0] rs1_l1,
    input  wire [ 4:0] rs2_l1,
    input  wire        ins_c_l1,
    input  wire        ins_lui_l1,
    input  wire        ins_auipc_l1,
    input  wire        ins_jal_l1,
    input  wire        ins_jalr_l1,
    input  wire        ins_beq_l1,
    input  wire        ins_bne_l1,
    input  wire        ins_blt_l1,
    input  wire        ins_bge_l1,
    input  wire        ins_bltu_l1,
    input  wire        ins_bgeu_l1,
    input  wire        ins_lb_l1,
    input  wire        ins_lh_l1,
    input  wire        ins_lw_l1,
    input  wire        ins_lbu_l1,
    input  wire        ins_lhu_l1,
    input  wire        ins_sb_l1,
    input  wire        ins_sh_l1,
    input  wire        ins_sw_l1,
    input  wire        ins_addi_l1,
    input  wire        ins_slti_l1,
    input  wire        ins_sltiu_l1,
    input  wire        ins_xori_l1,
    input  wire        ins_ori_l1,
    input  wire        ins_andi_l1,
    input  wire        ins_slli_l1,
    input  wire        ins_srli_l1,
    input  wire        ins_srai_l1,
    input  wire        ins_add_l1,
    input  wire        ins_sub_l1,
    input  wire        ins_sll_l1,
    input  wire        ins_slt_l1,
    input  wire        ins_sltu_l1,
    input  wire        ins_xor_l1,
    input  wire        ins_srl_l1,
    input  wire        ins_sra_l1,
    input  wire        ins_or_l1,
    input  wire        ins_and_l1,
    output reg  [31:0] pc_l2,
    output reg  [31:0] imm_l2,
    output reg  [ 4:0] rd_l2,
    output reg  [ 4:0] rs1_l2,
    output reg  [ 4:0] rs2_l2,
    output reg         ins_c_l2,
    output reg         ins_lui_l2,
    output reg         ins_auipc_l2,
    output reg         ins_jal_l2,
    output reg         ins_jalr_l2,
    output reg         ins_beq_l2,
    output reg         ins_bne_l2,
    output reg         ins_blt_l2,
    output reg         ins_bge_l2,
    output reg         ins_bltu_l2,
    output reg         ins_bgeu_l2,
    output reg         ins_lb_l2,
    output reg         ins_lh_l2,
    output reg         ins_lw_l2,
    output reg         ins_lbu_l2,
    output reg         ins_lhu_l2,
    output reg         ins_sb_l2,
    output reg         ins_sh_l2,
    output reg         ins_sw_l2,
    output reg         ins_addi_l2,
    output reg         ins_slti_l2,
    output reg         ins_sltiu_l2,
    output reg         ins_xori_l2,
    output reg         ins_ori_l2,
    output reg         ins_andi_l2,
    output reg         ins_slli_l2,
    output reg         ins_srli_l2,
    output reg         ins_srai_l2,
    output reg         ins_add_l2,
    output reg         ins_sub_l2,
    output reg         ins_sll_l2,
    output reg         ins_slt_l2,
    output reg         ins_sltu_l2,
    output reg         ins_xor_l2,
    output reg         ins_srl_l2,
    output reg         ins_sra_l2,
    output reg         ins_or_l2,
    output reg         ins_and_l2
);

endmodule
